`ifndef INC_UVM_INC
`define INC_UVM_INC

import uvm_pkg::*;

`include "test_pkg.sv"

import test_pkg::*;

`endif