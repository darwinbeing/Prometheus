`ifndef INC_TEST_PKG
`define INC_TEST_PKG

`include "env_pkg.sv"

package test_pkg;
	import uvm_pkg::*;

endpackage



`endif